//
// Template for UVM-compliant testcase

`ifndef TEST__SV
`define TEST__SV

typedef class top_env_env;

class top_env_test extends uvm_test;

  `uvm_component_utils(top_env_test)

  top_env_env env;

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    env = top_env_env::type_id::create("env", this);
    uvm_config_db #(uvm_object_wrapper)::set(this, "env.master_agent.mast_sqr.run_phase",
                    "default_sequence", my_mst_sequencer_sequence_library::get_type()); 
  endfunction

endclass : top_env_test

`endif //TEST__SV

